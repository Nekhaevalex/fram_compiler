
* cell 
* pin new_pin
.SUBCKT  2
* net 1 new_net
* device instance name r0 *1 0,0 pmos25
XD_name pmos25 PARAMS:
.ENDS 
