* Declare basic devices
* Memory cell subcuircuit
.SUBCKT memory_cell bl wl pl gnd
MM0 net6 wn bl gnd nsvt25 w=0.4 l=0.28
*X0 pl net6 conder Ec=1.9 dT=1e-09 l=5e-07 w=5e-07 p00=0.25
.ENDS memory_cell

* sense_amp subcuircuit
.SUBCKT sense_amp in ref seb nb nt vdd gnd
M3 nb seb gnd gnd nsvt25 w=0.4 l=0.28
M2 gnd seb nt gnd nsvt25 w=0.4 l=0.28
M1 nt nb gnd gnd nsvt25 w=0.4 l=0.28
M0 gnd nt nb gnd nsvt25 w=0.4 l=0.28
M8 net25 seb vdd vdd psvt25 w=0.4 l=0.28
M7 net25 ref net33 vdd psvt25 w=0.4 l=0.28
M6 net29 in net25 vdd psvt25 w=0.4 l=0.28
M5 nt nb net33 vdd psvt25 w=0.4 l=0.28
M4 net29 nt nb vdd psvt25 w=0.4 l=0.28
* SA
.ENDS
* Library name: fram_cells3
* Cell name: top_driver
* View name: schematic
.SUBCKT top_driver out in bl_gnd vdd gnd
M0 out in vdd vdd psvt25 w=2.0 l=0.28
M3 out in net19 gnd nsvt25 w=2.0 l=0.28
M1 net19 bl_gnd gnd gnd nsvt25 w=2.0 l=0.28
.ENDS top_driver// Generated for: spectre
// Generated on: Apr 23 22:43:59 2020
// Design library name: fram_cells5
// Design cell name: mos_pair_t
// Design view name: schematic

// Library name: fram_cells5
// Cell name: mos_pair
// View name: schematic
subckt mos_pair gnd in out_n out_p vdd
M0 (out_n in gnd gnd) nsvt25 w=0.4 l=0.28
M1 (out_p in vdd vdd) psvt25 w=0.4 l=0.28
ends mos_pair
// End of subcircuit definition.

// Library name: fram_cells5
// Cell name: mos_pair_t
// View name: schematic* Declare subcurcuits
* Declare instances
X0 bl0 wl0 pl0 gnd memory_cell
X1 bl0 wl1 pl1 gnd memory_cell
X2 bl0 wl2 pl2 gnd memory_cell
X3 bl0 wl3 pl3 gnd memory_cell
X4 bl0 wl4 pl4 gnd memory_cell
X5 bl0 wl5 pl5 gnd memory_cell
X6 bl0 wl6 pl6 gnd memory_cell
X7 bl0 wl7 pl7 gnd memory_cell
X8 bl0 wl8 pl8 gnd memory_cell
X9 bl0 wl9 pl9 gnd memory_cell
X10 bl0 wl10 pl10 gnd memory_cell
X11 bl0 wl11 pl11 gnd memory_cell
X12 bl0 wl12 pl12 gnd memory_cell
X13 bl0 wl13 pl13 gnd memory_cell
X14 bl0 wl14 pl14 gnd memory_cell
X15 bl0 wl15 pl15 gnd memory_cell
X16 bl0 wl16 pl16 gnd memory_cell
X17 bl0 wl17 pl17 gnd memory_cell
X18 bl0 wl18 pl18 gnd memory_cell
X19 bl0 wl19 pl19 gnd memory_cell
X20 bl0 wl20 pl20 gnd memory_cell
X21 bl0 wl21 pl21 gnd memory_cell
X22 bl0 wl22 pl22 gnd memory_cell
X23 bl0 wl23 pl23 gnd memory_cell
X24 bl0 wl24 pl24 gnd memory_cell
X25 bl0 wl25 pl25 gnd memory_cell
X26 bl0 wl26 pl26 gnd memory_cell
X27 bl0 wl27 pl27 gnd memory_cell
X28 bl0 wl28 pl28 gnd memory_cell
X29 bl0 wl29 pl29 gnd memory_cell
X30 bl0 wl30 pl30 gnd memory_cell
X31 bl0 wl31 pl31 gnd memory_cell
X32 bl1 wl0 pl0 gnd memory_cell
X33 bl1 wl1 pl1 gnd memory_cell
X34 bl1 wl2 pl2 gnd memory_cell
X35 bl1 wl3 pl3 gnd memory_cell
X36 bl1 wl4 pl4 gnd memory_cell
X37 bl1 wl5 pl5 gnd memory_cell
X38 bl1 wl6 pl6 gnd memory_cell
X39 bl1 wl7 pl7 gnd memory_cell
X40 bl1 wl8 pl8 gnd memory_cell
X41 bl1 wl9 pl9 gnd memory_cell
X42 bl1 wl10 pl10 gnd memory_cell
X43 bl1 wl11 pl11 gnd memory_cell
X44 bl1 wl12 pl12 gnd memory_cell
X45 bl1 wl13 pl13 gnd memory_cell
X46 bl1 wl14 pl14 gnd memory_cell
X47 bl1 wl15 pl15 gnd memory_cell
X48 bl1 wl16 pl16 gnd memory_cell
X49 bl1 wl17 pl17 gnd memory_cell
X50 bl1 wl18 pl18 gnd memory_cell
X51 bl1 wl19 pl19 gnd memory_cell
X52 bl1 wl20 pl20 gnd memory_cell
X53 bl1 wl21 pl21 gnd memory_cell
X54 bl1 wl22 pl22 gnd memory_cell
X55 bl1 wl23 pl23 gnd memory_cell
X56 bl1 wl24 pl24 gnd memory_cell
X57 bl1 wl25 pl25 gnd memory_cell
X58 bl1 wl26 pl26 gnd memory_cell
X59 bl1 wl27 pl27 gnd memory_cell
X60 bl1 wl28 pl28 gnd memory_cell
X61 bl1 wl29 pl29 gnd memory_cell
X62 bl1 wl30 pl30 gnd memory_cell
X63 bl1 wl31 pl31 gnd memory_cell
X64 bl2 wl0 pl0 gnd memory_cell
X65 bl2 wl1 pl1 gnd memory_cell
X66 bl2 wl2 pl2 gnd memory_cell
X67 bl2 wl3 pl3 gnd memory_cell
X68 bl2 wl4 pl4 gnd memory_cell
X69 bl2 wl5 pl5 gnd memory_cell
X70 bl2 wl6 pl6 gnd memory_cell
X71 bl2 wl7 pl7 gnd memory_cell
X72 bl2 wl8 pl8 gnd memory_cell
X73 bl2 wl9 pl9 gnd memory_cell
X74 bl2 wl10 pl10 gnd memory_cell
X75 bl2 wl11 pl11 gnd memory_cell
X76 bl2 wl12 pl12 gnd memory_cell
X77 bl2 wl13 pl13 gnd memory_cell
X78 bl2 wl14 pl14 gnd memory_cell
X79 bl2 wl15 pl15 gnd memory_cell
X80 bl2 wl16 pl16 gnd memory_cell
X81 bl2 wl17 pl17 gnd memory_cell
X82 bl2 wl18 pl18 gnd memory_cell
X83 bl2 wl19 pl19 gnd memory_cell
X84 bl2 wl20 pl20 gnd memory_cell
X85 bl2 wl21 pl21 gnd memory_cell
X86 bl2 wl22 pl22 gnd memory_cell
X87 bl2 wl23 pl23 gnd memory_cell
X88 bl2 wl24 pl24 gnd memory_cell
X89 bl2 wl25 pl25 gnd memory_cell
X90 bl2 wl26 pl26 gnd memory_cell
X91 bl2 wl27 pl27 gnd memory_cell
X92 bl2 wl28 pl28 gnd memory_cell
X93 bl2 wl29 pl29 gnd memory_cell
X94 bl2 wl30 pl30 gnd memory_cell
X95 bl2 wl31 pl31 gnd memory_cell
X96 bl3 wl0 pl0 gnd memory_cell
X97 bl3 wl1 pl1 gnd memory_cell
X98 bl3 wl2 pl2 gnd memory_cell
X99 bl3 wl3 pl3 gnd memory_cell
X100 bl3 wl4 pl4 gnd memory_cell
X101 bl3 wl5 pl5 gnd memory_cell
X102 bl3 wl6 pl6 gnd memory_cell
X103 bl3 wl7 pl7 gnd memory_cell
X104 bl3 wl8 pl8 gnd memory_cell
X105 bl3 wl9 pl9 gnd memory_cell
X106 bl3 wl10 pl10 gnd memory_cell
X107 bl3 wl11 pl11 gnd memory_cell
X108 bl3 wl12 pl12 gnd memory_cell
X109 bl3 wl13 pl13 gnd memory_cell
X110 bl3 wl14 pl14 gnd memory_cell
X111 bl3 wl15 pl15 gnd memory_cell
X112 bl3 wl16 pl16 gnd memory_cell
X113 bl3 wl17 pl17 gnd memory_cell
X114 bl3 wl18 pl18 gnd memory_cell
X115 bl3 wl19 pl19 gnd memory_cell
X116 bl3 wl20 pl20 gnd memory_cell
X117 bl3 wl21 pl21 gnd memory_cell
X118 bl3 wl22 pl22 gnd memory_cell
X119 bl3 wl23 pl23 gnd memory_cell
X120 bl3 wl24 pl24 gnd memory_cell
X121 bl3 wl25 pl25 gnd memory_cell
X122 bl3 wl26 pl26 gnd memory_cell
X123 bl3 wl27 pl27 gnd memory_cell
X124 bl3 wl28 pl28 gnd memory_cell
X125 bl3 wl29 pl29 gnd memory_cell
X126 bl3 wl30 pl30 gnd memory_cell
X127 bl3 wl31 pl31 gnd memory_cell
X128 bl4 wl0 pl0 gnd memory_cell
X129 bl4 wl1 pl1 gnd memory_cell
X130 bl4 wl2 pl2 gnd memory_cell
X131 bl4 wl3 pl3 gnd memory_cell
X132 bl4 wl4 pl4 gnd memory_cell
X133 bl4 wl5 pl5 gnd memory_cell
X134 bl4 wl6 pl6 gnd memory_cell
X135 bl4 wl7 pl7 gnd memory_cell
X136 bl4 wl8 pl8 gnd memory_cell
X137 bl4 wl9 pl9 gnd memory_cell
X138 bl4 wl10 pl10 gnd memory_cell
X139 bl4 wl11 pl11 gnd memory_cell
X140 bl4 wl12 pl12 gnd memory_cell
X141 bl4 wl13 pl13 gnd memory_cell
X142 bl4 wl14 pl14 gnd memory_cell
X143 bl4 wl15 pl15 gnd memory_cell
X144 bl4 wl16 pl16 gnd memory_cell
X145 bl4 wl17 pl17 gnd memory_cell
X146 bl4 wl18 pl18 gnd memory_cell
X147 bl4 wl19 pl19 gnd memory_cell
X148 bl4 wl20 pl20 gnd memory_cell
X149 bl4 wl21 pl21 gnd memory_cell
X150 bl4 wl22 pl22 gnd memory_cell
X151 bl4 wl23 pl23 gnd memory_cell
X152 bl4 wl24 pl24 gnd memory_cell
X153 bl4 wl25 pl25 gnd memory_cell
X154 bl4 wl26 pl26 gnd memory_cell
X155 bl4 wl27 pl27 gnd memory_cell
X156 bl4 wl28 pl28 gnd memory_cell
X157 bl4 wl29 pl29 gnd memory_cell
X158 bl4 wl30 pl30 gnd memory_cell
X159 bl4 wl31 pl31 gnd memory_cell
X160 bl5 wl0 pl0 gnd memory_cell
X161 bl5 wl1 pl1 gnd memory_cell
X162 bl5 wl2 pl2 gnd memory_cell
X163 bl5 wl3 pl3 gnd memory_cell
X164 bl5 wl4 pl4 gnd memory_cell
X165 bl5 wl5 pl5 gnd memory_cell
X166 bl5 wl6 pl6 gnd memory_cell
X167 bl5 wl7 pl7 gnd memory_cell
X168 bl5 wl8 pl8 gnd memory_cell
X169 bl5 wl9 pl9 gnd memory_cell
X170 bl5 wl10 pl10 gnd memory_cell
X171 bl5 wl11 pl11 gnd memory_cell
X172 bl5 wl12 pl12 gnd memory_cell
X173 bl5 wl13 pl13 gnd memory_cell
X174 bl5 wl14 pl14 gnd memory_cell
X175 bl5 wl15 pl15 gnd memory_cell
X176 bl5 wl16 pl16 gnd memory_cell
X177 bl5 wl17 pl17 gnd memory_cell
X178 bl5 wl18 pl18 gnd memory_cell
X179 bl5 wl19 pl19 gnd memory_cell
X180 bl5 wl20 pl20 gnd memory_cell
X181 bl5 wl21 pl21 gnd memory_cell
X182 bl5 wl22 pl22 gnd memory_cell
X183 bl5 wl23 pl23 gnd memory_cell
X184 bl5 wl24 pl24 gnd memory_cell
X185 bl5 wl25 pl25 gnd memory_cell
X186 bl5 wl26 pl26 gnd memory_cell
X187 bl5 wl27 pl27 gnd memory_cell
X188 bl5 wl28 pl28 gnd memory_cell
X189 bl5 wl29 pl29 gnd memory_cell
X190 bl5 wl30 pl30 gnd memory_cell
X191 bl5 wl31 pl31 gnd memory_cell
X192 bl6 wl0 pl0 gnd memory_cell
X193 bl6 wl1 pl1 gnd memory_cell
X194 bl6 wl2 pl2 gnd memory_cell
X195 bl6 wl3 pl3 gnd memory_cell
X196 bl6 wl4 pl4 gnd memory_cell
X197 bl6 wl5 pl5 gnd memory_cell
X198 bl6 wl6 pl6 gnd memory_cell
X199 bl6 wl7 pl7 gnd memory_cell
X200 bl6 wl8 pl8 gnd memory_cell
X201 bl6 wl9 pl9 gnd memory_cell
X202 bl6 wl10 pl10 gnd memory_cell
X203 bl6 wl11 pl11 gnd memory_cell
X204 bl6 wl12 pl12 gnd memory_cell
X205 bl6 wl13 pl13 gnd memory_cell
X206 bl6 wl14 pl14 gnd memory_cell
X207 bl6 wl15 pl15 gnd memory_cell
X208 bl6 wl16 pl16 gnd memory_cell
X209 bl6 wl17 pl17 gnd memory_cell
X210 bl6 wl18 pl18 gnd memory_cell
X211 bl6 wl19 pl19 gnd memory_cell
X212 bl6 wl20 pl20 gnd memory_cell
X213 bl6 wl21 pl21 gnd memory_cell
X214 bl6 wl22 pl22 gnd memory_cell
X215 bl6 wl23 pl23 gnd memory_cell
X216 bl6 wl24 pl24 gnd memory_cell
X217 bl6 wl25 pl25 gnd memory_cell
X218 bl6 wl26 pl26 gnd memory_cell
X219 bl6 wl27 pl27 gnd memory_cell
X220 bl6 wl28 pl28 gnd memory_cell
X221 bl6 wl29 pl29 gnd memory_cell
X222 bl6 wl30 pl30 gnd memory_cell
X223 bl6 wl31 pl31 gnd memory_cell
X224 bl7 wl0 pl0 gnd memory_cell
X225 bl7 wl1 pl1 gnd memory_cell
X226 bl7 wl2 pl2 gnd memory_cell
X227 bl7 wl3 pl3 gnd memory_cell
X228 bl7 wl4 pl4 gnd memory_cell
X229 bl7 wl5 pl5 gnd memory_cell
X230 bl7 wl6 pl6 gnd memory_cell
X231 bl7 wl7 pl7 gnd memory_cell
X232 bl7 wl8 pl8 gnd memory_cell
X233 bl7 wl9 pl9 gnd memory_cell
X234 bl7 wl10 pl10 gnd memory_cell
X235 bl7 wl11 pl11 gnd memory_cell
X236 bl7 wl12 pl12 gnd memory_cell
X237 bl7 wl13 pl13 gnd memory_cell
X238 bl7 wl14 pl14 gnd memory_cell
X239 bl7 wl15 pl15 gnd memory_cell
X240 bl7 wl16 pl16 gnd memory_cell
X241 bl7 wl17 pl17 gnd memory_cell
X242 bl7 wl18 pl18 gnd memory_cell
X243 bl7 wl19 pl19 gnd memory_cell
X244 bl7 wl20 pl20 gnd memory_cell
X245 bl7 wl21 pl21 gnd memory_cell
X246 bl7 wl22 pl22 gnd memory_cell
X247 bl7 wl23 pl23 gnd memory_cell
X248 bl7 wl24 pl24 gnd memory_cell
X249 bl7 wl25 pl25 gnd memory_cell
X250 bl7 wl26 pl26 gnd memory_cell
X251 bl7 wl27 pl27 gnd memory_cell
X252 bl7 wl28 pl28 gnd memory_cell
X253 bl7 wl29 pl29 gnd memory_cell
X254 bl7 wl30 pl30 gnd memory_cell
X255 bl7 wl31 pl31 gnd memory_cell
X256 bl8 wl0 pl0 gnd memory_cell
X257 bl8 wl1 pl1 gnd memory_cell
X258 bl8 wl2 pl2 gnd memory_cell
X259 bl8 wl3 pl3 gnd memory_cell
X260 bl8 wl4 pl4 gnd memory_cell
X261 bl8 wl5 pl5 gnd memory_cell
X262 bl8 wl6 pl6 gnd memory_cell
X263 bl8 wl7 pl7 gnd memory_cell
X264 bl8 wl8 pl8 gnd memory_cell
X265 bl8 wl9 pl9 gnd memory_cell
X266 bl8 wl10 pl10 gnd memory_cell
X267 bl8 wl11 pl11 gnd memory_cell
X268 bl8 wl12 pl12 gnd memory_cell
X269 bl8 wl13 pl13 gnd memory_cell
X270 bl8 wl14 pl14 gnd memory_cell
X271 bl8 wl15 pl15 gnd memory_cell
X272 bl8 wl16 pl16 gnd memory_cell
X273 bl8 wl17 pl17 gnd memory_cell
X274 bl8 wl18 pl18 gnd memory_cell
X275 bl8 wl19 pl19 gnd memory_cell
X276 bl8 wl20 pl20 gnd memory_cell
X277 bl8 wl21 pl21 gnd memory_cell
X278 bl8 wl22 pl22 gnd memory_cell
X279 bl8 wl23 pl23 gnd memory_cell
X280 bl8 wl24 pl24 gnd memory_cell
X281 bl8 wl25 pl25 gnd memory_cell
X282 bl8 wl26 pl26 gnd memory_cell
X283 bl8 wl27 pl27 gnd memory_cell
X284 bl8 wl28 pl28 gnd memory_cell
X285 bl8 wl29 pl29 gnd memory_cell
X286 bl8 wl30 pl30 gnd memory_cell
X287 bl8 wl31 pl31 gnd memory_cell
X288 bl9 wl0 pl0 gnd memory_cell
X289 bl9 wl1 pl1 gnd memory_cell
X290 bl9 wl2 pl2 gnd memory_cell
X291 bl9 wl3 pl3 gnd memory_cell
X292 bl9 wl4 pl4 gnd memory_cell
X293 bl9 wl5 pl5 gnd memory_cell
X294 bl9 wl6 pl6 gnd memory_cell
X295 bl9 wl7 pl7 gnd memory_cell
X296 bl9 wl8 pl8 gnd memory_cell
X297 bl9 wl9 pl9 gnd memory_cell
X298 bl9 wl10 pl10 gnd memory_cell
X299 bl9 wl11 pl11 gnd memory_cell
X300 bl9 wl12 pl12 gnd memory_cell
X301 bl9 wl13 pl13 gnd memory_cell
X302 bl9 wl14 pl14 gnd memory_cell
X303 bl9 wl15 pl15 gnd memory_cell
X304 bl9 wl16 pl16 gnd memory_cell
X305 bl9 wl17 pl17 gnd memory_cell
X306 bl9 wl18 pl18 gnd memory_cell
X307 bl9 wl19 pl19 gnd memory_cell
X308 bl9 wl20 pl20 gnd memory_cell
X309 bl9 wl21 pl21 gnd memory_cell
X310 bl9 wl22 pl22 gnd memory_cell
X311 bl9 wl23 pl23 gnd memory_cell
X312 bl9 wl24 pl24 gnd memory_cell
X313 bl9 wl25 pl25 gnd memory_cell
X314 bl9 wl26 pl26 gnd memory_cell
X315 bl9 wl27 pl27 gnd memory_cell
X316 bl9 wl28 pl28 gnd memory_cell
X317 bl9 wl29 pl29 gnd memory_cell
X318 bl9 wl30 pl30 gnd memory_cell
X319 bl9 wl31 pl31 gnd memory_cell
X320 bl10 wl0 pl0 gnd memory_cell
X321 bl10 wl1 pl1 gnd memory_cell
X322 bl10 wl2 pl2 gnd memory_cell
X323 bl10 wl3 pl3 gnd memory_cell
X324 bl10 wl4 pl4 gnd memory_cell
X325 bl10 wl5 pl5 gnd memory_cell
X326 bl10 wl6 pl6 gnd memory_cell
X327 bl10 wl7 pl7 gnd memory_cell
X328 bl10 wl8 pl8 gnd memory_cell
X329 bl10 wl9 pl9 gnd memory_cell
X330 bl10 wl10 pl10 gnd memory_cell
X331 bl10 wl11 pl11 gnd memory_cell
X332 bl10 wl12 pl12 gnd memory_cell
X333 bl10 wl13 pl13 gnd memory_cell
X334 bl10 wl14 pl14 gnd memory_cell
X335 bl10 wl15 pl15 gnd memory_cell
X336 bl10 wl16 pl16 gnd memory_cell
X337 bl10 wl17 pl17 gnd memory_cell
X338 bl10 wl18 pl18 gnd memory_cell
X339 bl10 wl19 pl19 gnd memory_cell
X340 bl10 wl20 pl20 gnd memory_cell
X341 bl10 wl21 pl21 gnd memory_cell
X342 bl10 wl22 pl22 gnd memory_cell
X343 bl10 wl23 pl23 gnd memory_cell
X344 bl10 wl24 pl24 gnd memory_cell
X345 bl10 wl25 pl25 gnd memory_cell
X346 bl10 wl26 pl26 gnd memory_cell
X347 bl10 wl27 pl27 gnd memory_cell
X348 bl10 wl28 pl28 gnd memory_cell
X349 bl10 wl29 pl29 gnd memory_cell
X350 bl10 wl30 pl30 gnd memory_cell
X351 bl10 wl31 pl31 gnd memory_cell
X352 bl11 wl0 pl0 gnd memory_cell
X353 bl11 wl1 pl1 gnd memory_cell
X354 bl11 wl2 pl2 gnd memory_cell
X355 bl11 wl3 pl3 gnd memory_cell
X356 bl11 wl4 pl4 gnd memory_cell
X357 bl11 wl5 pl5 gnd memory_cell
X358 bl11 wl6 pl6 gnd memory_cell
X359 bl11 wl7 pl7 gnd memory_cell
X360 bl11 wl8 pl8 gnd memory_cell
X361 bl11 wl9 pl9 gnd memory_cell
X362 bl11 wl10 pl10 gnd memory_cell
X363 bl11 wl11 pl11 gnd memory_cell
X364 bl11 wl12 pl12 gnd memory_cell
X365 bl11 wl13 pl13 gnd memory_cell
X366 bl11 wl14 pl14 gnd memory_cell
X367 bl11 wl15 pl15 gnd memory_cell
X368 bl11 wl16 pl16 gnd memory_cell
X369 bl11 wl17 pl17 gnd memory_cell
X370 bl11 wl18 pl18 gnd memory_cell
X371 bl11 wl19 pl19 gnd memory_cell
X372 bl11 wl20 pl20 gnd memory_cell
X373 bl11 wl21 pl21 gnd memory_cell
X374 bl11 wl22 pl22 gnd memory_cell
X375 bl11 wl23 pl23 gnd memory_cell
X376 bl11 wl24 pl24 gnd memory_cell
X377 bl11 wl25 pl25 gnd memory_cell
X378 bl11 wl26 pl26 gnd memory_cell
X379 bl11 wl27 pl27 gnd memory_cell
X380 bl11 wl28 pl28 gnd memory_cell
X381 bl11 wl29 pl29 gnd memory_cell
X382 bl11 wl30 pl30 gnd memory_cell
X383 bl11 wl31 pl31 gnd memory_cell
X384 bl12 wl0 pl0 gnd memory_cell
X385 bl12 wl1 pl1 gnd memory_cell
X386 bl12 wl2 pl2 gnd memory_cell
X387 bl12 wl3 pl3 gnd memory_cell
X388 bl12 wl4 pl4 gnd memory_cell
X389 bl12 wl5 pl5 gnd memory_cell
X390 bl12 wl6 pl6 gnd memory_cell
X391 bl12 wl7 pl7 gnd memory_cell
X392 bl12 wl8 pl8 gnd memory_cell
X393 bl12 wl9 pl9 gnd memory_cell
X394 bl12 wl10 pl10 gnd memory_cell
X395 bl12 wl11 pl11 gnd memory_cell
X396 bl12 wl12 pl12 gnd memory_cell
X397 bl12 wl13 pl13 gnd memory_cell
X398 bl12 wl14 pl14 gnd memory_cell
X399 bl12 wl15 pl15 gnd memory_cell
X400 bl12 wl16 pl16 gnd memory_cell
X401 bl12 wl17 pl17 gnd memory_cell
X402 bl12 wl18 pl18 gnd memory_cell
X403 bl12 wl19 pl19 gnd memory_cell
X404 bl12 wl20 pl20 gnd memory_cell
X405 bl12 wl21 pl21 gnd memory_cell
X406 bl12 wl22 pl22 gnd memory_cell
X407 bl12 wl23 pl23 gnd memory_cell
X408 bl12 wl24 pl24 gnd memory_cell
X409 bl12 wl25 pl25 gnd memory_cell
X410 bl12 wl26 pl26 gnd memory_cell
X411 bl12 wl27 pl27 gnd memory_cell
X412 bl12 wl28 pl28 gnd memory_cell
X413 bl12 wl29 pl29 gnd memory_cell
X414 bl12 wl30 pl30 gnd memory_cell
X415 bl12 wl31 pl31 gnd memory_cell
X416 bl13 wl0 pl0 gnd memory_cell
X417 bl13 wl1 pl1 gnd memory_cell
X418 bl13 wl2 pl2 gnd memory_cell
X419 bl13 wl3 pl3 gnd memory_cell
X420 bl13 wl4 pl4 gnd memory_cell
X421 bl13 wl5 pl5 gnd memory_cell
X422 bl13 wl6 pl6 gnd memory_cell
X423 bl13 wl7 pl7 gnd memory_cell
X424 bl13 wl8 pl8 gnd memory_cell
X425 bl13 wl9 pl9 gnd memory_cell
X426 bl13 wl10 pl10 gnd memory_cell
X427 bl13 wl11 pl11 gnd memory_cell
X428 bl13 wl12 pl12 gnd memory_cell
X429 bl13 wl13 pl13 gnd memory_cell
X430 bl13 wl14 pl14 gnd memory_cell
X431 bl13 wl15 pl15 gnd memory_cell
X432 bl13 wl16 pl16 gnd memory_cell
X433 bl13 wl17 pl17 gnd memory_cell
X434 bl13 wl18 pl18 gnd memory_cell
X435 bl13 wl19 pl19 gnd memory_cell
X436 bl13 wl20 pl20 gnd memory_cell
X437 bl13 wl21 pl21 gnd memory_cell
X438 bl13 wl22 pl22 gnd memory_cell
X439 bl13 wl23 pl23 gnd memory_cell
X440 bl13 wl24 pl24 gnd memory_cell
X441 bl13 wl25 pl25 gnd memory_cell
X442 bl13 wl26 pl26 gnd memory_cell
X443 bl13 wl27 pl27 gnd memory_cell
X444 bl13 wl28 pl28 gnd memory_cell
X445 bl13 wl29 pl29 gnd memory_cell
X446 bl13 wl30 pl30 gnd memory_cell
X447 bl13 wl31 pl31 gnd memory_cell
X448 bl14 wl0 pl0 gnd memory_cell
X449 bl14 wl1 pl1 gnd memory_cell
X450 bl14 wl2 pl2 gnd memory_cell
X451 bl14 wl3 pl3 gnd memory_cell
X452 bl14 wl4 pl4 gnd memory_cell
X453 bl14 wl5 pl5 gnd memory_cell
X454 bl14 wl6 pl6 gnd memory_cell
X455 bl14 wl7 pl7 gnd memory_cell
X456 bl14 wl8 pl8 gnd memory_cell
X457 bl14 wl9 pl9 gnd memory_cell
X458 bl14 wl10 pl10 gnd memory_cell
X459 bl14 wl11 pl11 gnd memory_cell
X460 bl14 wl12 pl12 gnd memory_cell
X461 bl14 wl13 pl13 gnd memory_cell
X462 bl14 wl14 pl14 gnd memory_cell
X463 bl14 wl15 pl15 gnd memory_cell
X464 bl14 wl16 pl16 gnd memory_cell
X465 bl14 wl17 pl17 gnd memory_cell
X466 bl14 wl18 pl18 gnd memory_cell
X467 bl14 wl19 pl19 gnd memory_cell
X468 bl14 wl20 pl20 gnd memory_cell
X469 bl14 wl21 pl21 gnd memory_cell
X470 bl14 wl22 pl22 gnd memory_cell
X471 bl14 wl23 pl23 gnd memory_cell
X472 bl14 wl24 pl24 gnd memory_cell
X473 bl14 wl25 pl25 gnd memory_cell
X474 bl14 wl26 pl26 gnd memory_cell
X475 bl14 wl27 pl27 gnd memory_cell
X476 bl14 wl28 pl28 gnd memory_cell
X477 bl14 wl29 pl29 gnd memory_cell
X478 bl14 wl30 pl30 gnd memory_cell
X479 bl14 wl31 pl31 gnd memory_cell
X480 bl15 wl0 pl0 gnd memory_cell
X481 bl15 wl1 pl1 gnd memory_cell
X482 bl15 wl2 pl2 gnd memory_cell
X483 bl15 wl3 pl3 gnd memory_cell
X484 bl15 wl4 pl4 gnd memory_cell
X485 bl15 wl5 pl5 gnd memory_cell
X486 bl15 wl6 pl6 gnd memory_cell
X487 bl15 wl7 pl7 gnd memory_cell
X488 bl15 wl8 pl8 gnd memory_cell
X489 bl15 wl9 pl9 gnd memory_cell
X490 bl15 wl10 pl10 gnd memory_cell
X491 bl15 wl11 pl11 gnd memory_cell
X492 bl15 wl12 pl12 gnd memory_cell
X493 bl15 wl13 pl13 gnd memory_cell
X494 bl15 wl14 pl14 gnd memory_cell
X495 bl15 wl15 pl15 gnd memory_cell
X496 bl15 wl16 pl16 gnd memory_cell
X497 bl15 wl17 pl17 gnd memory_cell
X498 bl15 wl18 pl18 gnd memory_cell
X499 bl15 wl19 pl19 gnd memory_cell
X500 bl15 wl20 pl20 gnd memory_cell
X501 bl15 wl21 pl21 gnd memory_cell
X502 bl15 wl22 pl22 gnd memory_cell
X503 bl15 wl23 pl23 gnd memory_cell
X504 bl15 wl24 pl24 gnd memory_cell
X505 bl15 wl25 pl25 gnd memory_cell
X506 bl15 wl26 pl26 gnd memory_cell
X507 bl15 wl27 pl27 gnd memory_cell
X508 bl15 wl28 pl28 gnd memory_cell
X509 bl15 wl29 pl29 gnd memory_cell
X510 bl15 wl30 pl30 gnd memory_cell
X511 bl15 wl31 pl31 gnd memory_cell
X512 bl16 wl0 pl0 gnd memory_cell
X513 bl16 wl1 pl1 gnd memory_cell
X514 bl16 wl2 pl2 gnd memory_cell
X515 bl16 wl3 pl3 gnd memory_cell
X516 bl16 wl4 pl4 gnd memory_cell
X517 bl16 wl5 pl5 gnd memory_cell
X518 bl16 wl6 pl6 gnd memory_cell
X519 bl16 wl7 pl7 gnd memory_cell
X520 bl16 wl8 pl8 gnd memory_cell
X521 bl16 wl9 pl9 gnd memory_cell
X522 bl16 wl10 pl10 gnd memory_cell
X523 bl16 wl11 pl11 gnd memory_cell
X524 bl16 wl12 pl12 gnd memory_cell
X525 bl16 wl13 pl13 gnd memory_cell
X526 bl16 wl14 pl14 gnd memory_cell
X527 bl16 wl15 pl15 gnd memory_cell
X528 bl16 wl16 pl16 gnd memory_cell
X529 bl16 wl17 pl17 gnd memory_cell
X530 bl16 wl18 pl18 gnd memory_cell
X531 bl16 wl19 pl19 gnd memory_cell
X532 bl16 wl20 pl20 gnd memory_cell
X533 bl16 wl21 pl21 gnd memory_cell
X534 bl16 wl22 pl22 gnd memory_cell
X535 bl16 wl23 pl23 gnd memory_cell
X536 bl16 wl24 pl24 gnd memory_cell
X537 bl16 wl25 pl25 gnd memory_cell
X538 bl16 wl26 pl26 gnd memory_cell
X539 bl16 wl27 pl27 gnd memory_cell
X540 bl16 wl28 pl28 gnd memory_cell
X541 bl16 wl29 pl29 gnd memory_cell
X542 bl16 wl30 pl30 gnd memory_cell
X543 bl16 wl31 pl31 gnd memory_cell
X544 bl17 wl0 pl0 gnd memory_cell
X545 bl17 wl1 pl1 gnd memory_cell
X546 bl17 wl2 pl2 gnd memory_cell
X547 bl17 wl3 pl3 gnd memory_cell
X548 bl17 wl4 pl4 gnd memory_cell
X549 bl17 wl5 pl5 gnd memory_cell
X550 bl17 wl6 pl6 gnd memory_cell
X551 bl17 wl7 pl7 gnd memory_cell
X552 bl17 wl8 pl8 gnd memory_cell
X553 bl17 wl9 pl9 gnd memory_cell
X554 bl17 wl10 pl10 gnd memory_cell
X555 bl17 wl11 pl11 gnd memory_cell
X556 bl17 wl12 pl12 gnd memory_cell
X557 bl17 wl13 pl13 gnd memory_cell
X558 bl17 wl14 pl14 gnd memory_cell
X559 bl17 wl15 pl15 gnd memory_cell
X560 bl17 wl16 pl16 gnd memory_cell
X561 bl17 wl17 pl17 gnd memory_cell
X562 bl17 wl18 pl18 gnd memory_cell
X563 bl17 wl19 pl19 gnd memory_cell
X564 bl17 wl20 pl20 gnd memory_cell
X565 bl17 wl21 pl21 gnd memory_cell
X566 bl17 wl22 pl22 gnd memory_cell
X567 bl17 wl23 pl23 gnd memory_cell
X568 bl17 wl24 pl24 gnd memory_cell
X569 bl17 wl25 pl25 gnd memory_cell
X570 bl17 wl26 pl26 gnd memory_cell
X571 bl17 wl27 pl27 gnd memory_cell
X572 bl17 wl28 pl28 gnd memory_cell
X573 bl17 wl29 pl29 gnd memory_cell
X574 bl17 wl30 pl30 gnd memory_cell
X575 bl17 wl31 pl31 gnd memory_cell
X576 bl18 wl0 pl0 gnd memory_cell
X577 bl18 wl1 pl1 gnd memory_cell
X578 bl18 wl2 pl2 gnd memory_cell
X579 bl18 wl3 pl3 gnd memory_cell
X580 bl18 wl4 pl4 gnd memory_cell
X581 bl18 wl5 pl5 gnd memory_cell
X582 bl18 wl6 pl6 gnd memory_cell
X583 bl18 wl7 pl7 gnd memory_cell
X584 bl18 wl8 pl8 gnd memory_cell
X585 bl18 wl9 pl9 gnd memory_cell
X586 bl18 wl10 pl10 gnd memory_cell
X587 bl18 wl11 pl11 gnd memory_cell
X588 bl18 wl12 pl12 gnd memory_cell
X589 bl18 wl13 pl13 gnd memory_cell
X590 bl18 wl14 pl14 gnd memory_cell
X591 bl18 wl15 pl15 gnd memory_cell
X592 bl18 wl16 pl16 gnd memory_cell
X593 bl18 wl17 pl17 gnd memory_cell
X594 bl18 wl18 pl18 gnd memory_cell
X595 bl18 wl19 pl19 gnd memory_cell
X596 bl18 wl20 pl20 gnd memory_cell
X597 bl18 wl21 pl21 gnd memory_cell
X598 bl18 wl22 pl22 gnd memory_cell
X599 bl18 wl23 pl23 gnd memory_cell
X600 bl18 wl24 pl24 gnd memory_cell
X601 bl18 wl25 pl25 gnd memory_cell
X602 bl18 wl26 pl26 gnd memory_cell
X603 bl18 wl27 pl27 gnd memory_cell
X604 bl18 wl28 pl28 gnd memory_cell
X605 bl18 wl29 pl29 gnd memory_cell
X606 bl18 wl30 pl30 gnd memory_cell
X607 bl18 wl31 pl31 gnd memory_cell
X608 bl19 wl0 pl0 gnd memory_cell
X609 bl19 wl1 pl1 gnd memory_cell
X610 bl19 wl2 pl2 gnd memory_cell
X611 bl19 wl3 pl3 gnd memory_cell
X612 bl19 wl4 pl4 gnd memory_cell
X613 bl19 wl5 pl5 gnd memory_cell
X614 bl19 wl6 pl6 gnd memory_cell
X615 bl19 wl7 pl7 gnd memory_cell
X616 bl19 wl8 pl8 gnd memory_cell
X617 bl19 wl9 pl9 gnd memory_cell
X618 bl19 wl10 pl10 gnd memory_cell
X619 bl19 wl11 pl11 gnd memory_cell
X620 bl19 wl12 pl12 gnd memory_cell
X621 bl19 wl13 pl13 gnd memory_cell
X622 bl19 wl14 pl14 gnd memory_cell
X623 bl19 wl15 pl15 gnd memory_cell
X624 bl19 wl16 pl16 gnd memory_cell
X625 bl19 wl17 pl17 gnd memory_cell
X626 bl19 wl18 pl18 gnd memory_cell
X627 bl19 wl19 pl19 gnd memory_cell
X628 bl19 wl20 pl20 gnd memory_cell
X629 bl19 wl21 pl21 gnd memory_cell
X630 bl19 wl22 pl22 gnd memory_cell
X631 bl19 wl23 pl23 gnd memory_cell
X632 bl19 wl24 pl24 gnd memory_cell
X633 bl19 wl25 pl25 gnd memory_cell
X634 bl19 wl26 pl26 gnd memory_cell
X635 bl19 wl27 pl27 gnd memory_cell
X636 bl19 wl28 pl28 gnd memory_cell
X637 bl19 wl29 pl29 gnd memory_cell
X638 bl19 wl30 pl30 gnd memory_cell
X639 bl19 wl31 pl31 gnd memory_cell
X640 bl20 wl0 pl0 gnd memory_cell
X641 bl20 wl1 pl1 gnd memory_cell
X642 bl20 wl2 pl2 gnd memory_cell
X643 bl20 wl3 pl3 gnd memory_cell
X644 bl20 wl4 pl4 gnd memory_cell
X645 bl20 wl5 pl5 gnd memory_cell
X646 bl20 wl6 pl6 gnd memory_cell
X647 bl20 wl7 pl7 gnd memory_cell
X648 bl20 wl8 pl8 gnd memory_cell
X649 bl20 wl9 pl9 gnd memory_cell
X650 bl20 wl10 pl10 gnd memory_cell
X651 bl20 wl11 pl11 gnd memory_cell
X652 bl20 wl12 pl12 gnd memory_cell
X653 bl20 wl13 pl13 gnd memory_cell
X654 bl20 wl14 pl14 gnd memory_cell
X655 bl20 wl15 pl15 gnd memory_cell
X656 bl20 wl16 pl16 gnd memory_cell
X657 bl20 wl17 pl17 gnd memory_cell
X658 bl20 wl18 pl18 gnd memory_cell
X659 bl20 wl19 pl19 gnd memory_cell
X660 bl20 wl20 pl20 gnd memory_cell
X661 bl20 wl21 pl21 gnd memory_cell
X662 bl20 wl22 pl22 gnd memory_cell
X663 bl20 wl23 pl23 gnd memory_cell
X664 bl20 wl24 pl24 gnd memory_cell
X665 bl20 wl25 pl25 gnd memory_cell
X666 bl20 wl26 pl26 gnd memory_cell
X667 bl20 wl27 pl27 gnd memory_cell
X668 bl20 wl28 pl28 gnd memory_cell
X669 bl20 wl29 pl29 gnd memory_cell
X670 bl20 wl30 pl30 gnd memory_cell
X671 bl20 wl31 pl31 gnd memory_cell
X672 bl21 wl0 pl0 gnd memory_cell
X673 bl21 wl1 pl1 gnd memory_cell
X674 bl21 wl2 pl2 gnd memory_cell
X675 bl21 wl3 pl3 gnd memory_cell
X676 bl21 wl4 pl4 gnd memory_cell
X677 bl21 wl5 pl5 gnd memory_cell
X678 bl21 wl6 pl6 gnd memory_cell
X679 bl21 wl7 pl7 gnd memory_cell
X680 bl21 wl8 pl8 gnd memory_cell
X681 bl21 wl9 pl9 gnd memory_cell
X682 bl21 wl10 pl10 gnd memory_cell
X683 bl21 wl11 pl11 gnd memory_cell
X684 bl21 wl12 pl12 gnd memory_cell
X685 bl21 wl13 pl13 gnd memory_cell
X686 bl21 wl14 pl14 gnd memory_cell
X687 bl21 wl15 pl15 gnd memory_cell
X688 bl21 wl16 pl16 gnd memory_cell
X689 bl21 wl17 pl17 gnd memory_cell
X690 bl21 wl18 pl18 gnd memory_cell
X691 bl21 wl19 pl19 gnd memory_cell
X692 bl21 wl20 pl20 gnd memory_cell
X693 bl21 wl21 pl21 gnd memory_cell
X694 bl21 wl22 pl22 gnd memory_cell
X695 bl21 wl23 pl23 gnd memory_cell
X696 bl21 wl24 pl24 gnd memory_cell
X697 bl21 wl25 pl25 gnd memory_cell
X698 bl21 wl26 pl26 gnd memory_cell
X699 bl21 wl27 pl27 gnd memory_cell
X700 bl21 wl28 pl28 gnd memory_cell
X701 bl21 wl29 pl29 gnd memory_cell
X702 bl21 wl30 pl30 gnd memory_cell
X703 bl21 wl31 pl31 gnd memory_cell
X704 bl22 wl0 pl0 gnd memory_cell
X705 bl22 wl1 pl1 gnd memory_cell
X706 bl22 wl2 pl2 gnd memory_cell
X707 bl22 wl3 pl3 gnd memory_cell
X708 bl22 wl4 pl4 gnd memory_cell
X709 bl22 wl5 pl5 gnd memory_cell
X710 bl22 wl6 pl6 gnd memory_cell
X711 bl22 wl7 pl7 gnd memory_cell
X712 bl22 wl8 pl8 gnd memory_cell
X713 bl22 wl9 pl9 gnd memory_cell
X714 bl22 wl10 pl10 gnd memory_cell
X715 bl22 wl11 pl11 gnd memory_cell
X716 bl22 wl12 pl12 gnd memory_cell
X717 bl22 wl13 pl13 gnd memory_cell
X718 bl22 wl14 pl14 gnd memory_cell
X719 bl22 wl15 pl15 gnd memory_cell
X720 bl22 wl16 pl16 gnd memory_cell
X721 bl22 wl17 pl17 gnd memory_cell
X722 bl22 wl18 pl18 gnd memory_cell
X723 bl22 wl19 pl19 gnd memory_cell
X724 bl22 wl20 pl20 gnd memory_cell
X725 bl22 wl21 pl21 gnd memory_cell
X726 bl22 wl22 pl22 gnd memory_cell
X727 bl22 wl23 pl23 gnd memory_cell
X728 bl22 wl24 pl24 gnd memory_cell
X729 bl22 wl25 pl25 gnd memory_cell
X730 bl22 wl26 pl26 gnd memory_cell
X731 bl22 wl27 pl27 gnd memory_cell
X732 bl22 wl28 pl28 gnd memory_cell
X733 bl22 wl29 pl29 gnd memory_cell
X734 bl22 wl30 pl30 gnd memory_cell
X735 bl22 wl31 pl31 gnd memory_cell
X736 bl23 wl0 pl0 gnd memory_cell
X737 bl23 wl1 pl1 gnd memory_cell
X738 bl23 wl2 pl2 gnd memory_cell
X739 bl23 wl3 pl3 gnd memory_cell
X740 bl23 wl4 pl4 gnd memory_cell
X741 bl23 wl5 pl5 gnd memory_cell
X742 bl23 wl6 pl6 gnd memory_cell
X743 bl23 wl7 pl7 gnd memory_cell
X744 bl23 wl8 pl8 gnd memory_cell
X745 bl23 wl9 pl9 gnd memory_cell
X746 bl23 wl10 pl10 gnd memory_cell
X747 bl23 wl11 pl11 gnd memory_cell
X748 bl23 wl12 pl12 gnd memory_cell
X749 bl23 wl13 pl13 gnd memory_cell
X750 bl23 wl14 pl14 gnd memory_cell
X751 bl23 wl15 pl15 gnd memory_cell
X752 bl23 wl16 pl16 gnd memory_cell
X753 bl23 wl17 pl17 gnd memory_cell
X754 bl23 wl18 pl18 gnd memory_cell
X755 bl23 wl19 pl19 gnd memory_cell
X756 bl23 wl20 pl20 gnd memory_cell
X757 bl23 wl21 pl21 gnd memory_cell
X758 bl23 wl22 pl22 gnd memory_cell
X759 bl23 wl23 pl23 gnd memory_cell
X760 bl23 wl24 pl24 gnd memory_cell
X761 bl23 wl25 pl25 gnd memory_cell
X762 bl23 wl26 pl26 gnd memory_cell
X763 bl23 wl27 pl27 gnd memory_cell
X764 bl23 wl28 pl28 gnd memory_cell
X765 bl23 wl29 pl29 gnd memory_cell
X766 bl23 wl30 pl30 gnd memory_cell
X767 bl23 wl31 pl31 gnd memory_cell
X768 bl24 wl0 pl0 gnd memory_cell
X769 bl24 wl1 pl1 gnd memory_cell
X770 bl24 wl2 pl2 gnd memory_cell
X771 bl24 wl3 pl3 gnd memory_cell
X772 bl24 wl4 pl4 gnd memory_cell
X773 bl24 wl5 pl5 gnd memory_cell
X774 bl24 wl6 pl6 gnd memory_cell
X775 bl24 wl7 pl7 gnd memory_cell
X776 bl24 wl8 pl8 gnd memory_cell
X777 bl24 wl9 pl9 gnd memory_cell
X778 bl24 wl10 pl10 gnd memory_cell
X779 bl24 wl11 pl11 gnd memory_cell
X780 bl24 wl12 pl12 gnd memory_cell
X781 bl24 wl13 pl13 gnd memory_cell
X782 bl24 wl14 pl14 gnd memory_cell
X783 bl24 wl15 pl15 gnd memory_cell
X784 bl24 wl16 pl16 gnd memory_cell
X785 bl24 wl17 pl17 gnd memory_cell
X786 bl24 wl18 pl18 gnd memory_cell
X787 bl24 wl19 pl19 gnd memory_cell
X788 bl24 wl20 pl20 gnd memory_cell
X789 bl24 wl21 pl21 gnd memory_cell
X790 bl24 wl22 pl22 gnd memory_cell
X791 bl24 wl23 pl23 gnd memory_cell
X792 bl24 wl24 pl24 gnd memory_cell
X793 bl24 wl25 pl25 gnd memory_cell
X794 bl24 wl26 pl26 gnd memory_cell
X795 bl24 wl27 pl27 gnd memory_cell
X796 bl24 wl28 pl28 gnd memory_cell
X797 bl24 wl29 pl29 gnd memory_cell
X798 bl24 wl30 pl30 gnd memory_cell
X799 bl24 wl31 pl31 gnd memory_cell
X800 bl25 wl0 pl0 gnd memory_cell
X801 bl25 wl1 pl1 gnd memory_cell
X802 bl25 wl2 pl2 gnd memory_cell
X803 bl25 wl3 pl3 gnd memory_cell
X804 bl25 wl4 pl4 gnd memory_cell
X805 bl25 wl5 pl5 gnd memory_cell
X806 bl25 wl6 pl6 gnd memory_cell
X807 bl25 wl7 pl7 gnd memory_cell
X808 bl25 wl8 pl8 gnd memory_cell
X809 bl25 wl9 pl9 gnd memory_cell
X810 bl25 wl10 pl10 gnd memory_cell
X811 bl25 wl11 pl11 gnd memory_cell
X812 bl25 wl12 pl12 gnd memory_cell
X813 bl25 wl13 pl13 gnd memory_cell
X814 bl25 wl14 pl14 gnd memory_cell
X815 bl25 wl15 pl15 gnd memory_cell
X816 bl25 wl16 pl16 gnd memory_cell
X817 bl25 wl17 pl17 gnd memory_cell
X818 bl25 wl18 pl18 gnd memory_cell
X819 bl25 wl19 pl19 gnd memory_cell
X820 bl25 wl20 pl20 gnd memory_cell
X821 bl25 wl21 pl21 gnd memory_cell
X822 bl25 wl22 pl22 gnd memory_cell
X823 bl25 wl23 pl23 gnd memory_cell
X824 bl25 wl24 pl24 gnd memory_cell
X825 bl25 wl25 pl25 gnd memory_cell
X826 bl25 wl26 pl26 gnd memory_cell
X827 bl25 wl27 pl27 gnd memory_cell
X828 bl25 wl28 pl28 gnd memory_cell
X829 bl25 wl29 pl29 gnd memory_cell
X830 bl25 wl30 pl30 gnd memory_cell
X831 bl25 wl31 pl31 gnd memory_cell
X832 bl26 wl0 pl0 gnd memory_cell
X833 bl26 wl1 pl1 gnd memory_cell
X834 bl26 wl2 pl2 gnd memory_cell
X835 bl26 wl3 pl3 gnd memory_cell
X836 bl26 wl4 pl4 gnd memory_cell
X837 bl26 wl5 pl5 gnd memory_cell
X838 bl26 wl6 pl6 gnd memory_cell
X839 bl26 wl7 pl7 gnd memory_cell
X840 bl26 wl8 pl8 gnd memory_cell
X841 bl26 wl9 pl9 gnd memory_cell
X842 bl26 wl10 pl10 gnd memory_cell
X843 bl26 wl11 pl11 gnd memory_cell
X844 bl26 wl12 pl12 gnd memory_cell
X845 bl26 wl13 pl13 gnd memory_cell
X846 bl26 wl14 pl14 gnd memory_cell
X847 bl26 wl15 pl15 gnd memory_cell
X848 bl26 wl16 pl16 gnd memory_cell
X849 bl26 wl17 pl17 gnd memory_cell
X850 bl26 wl18 pl18 gnd memory_cell
X851 bl26 wl19 pl19 gnd memory_cell
X852 bl26 wl20 pl20 gnd memory_cell
X853 bl26 wl21 pl21 gnd memory_cell
X854 bl26 wl22 pl22 gnd memory_cell
X855 bl26 wl23 pl23 gnd memory_cell
X856 bl26 wl24 pl24 gnd memory_cell
X857 bl26 wl25 pl25 gnd memory_cell
X858 bl26 wl26 pl26 gnd memory_cell
X859 bl26 wl27 pl27 gnd memory_cell
X860 bl26 wl28 pl28 gnd memory_cell
X861 bl26 wl29 pl29 gnd memory_cell
X862 bl26 wl30 pl30 gnd memory_cell
X863 bl26 wl31 pl31 gnd memory_cell
X864 bl27 wl0 pl0 gnd memory_cell
X865 bl27 wl1 pl1 gnd memory_cell
X866 bl27 wl2 pl2 gnd memory_cell
X867 bl27 wl3 pl3 gnd memory_cell
X868 bl27 wl4 pl4 gnd memory_cell
X869 bl27 wl5 pl5 gnd memory_cell
X870 bl27 wl6 pl6 gnd memory_cell
X871 bl27 wl7 pl7 gnd memory_cell
X872 bl27 wl8 pl8 gnd memory_cell
X873 bl27 wl9 pl9 gnd memory_cell
X874 bl27 wl10 pl10 gnd memory_cell
X875 bl27 wl11 pl11 gnd memory_cell
X876 bl27 wl12 pl12 gnd memory_cell
X877 bl27 wl13 pl13 gnd memory_cell
X878 bl27 wl14 pl14 gnd memory_cell
X879 bl27 wl15 pl15 gnd memory_cell
X880 bl27 wl16 pl16 gnd memory_cell
X881 bl27 wl17 pl17 gnd memory_cell
X882 bl27 wl18 pl18 gnd memory_cell
X883 bl27 wl19 pl19 gnd memory_cell
X884 bl27 wl20 pl20 gnd memory_cell
X885 bl27 wl21 pl21 gnd memory_cell
X886 bl27 wl22 pl22 gnd memory_cell
X887 bl27 wl23 pl23 gnd memory_cell
X888 bl27 wl24 pl24 gnd memory_cell
X889 bl27 wl25 pl25 gnd memory_cell
X890 bl27 wl26 pl26 gnd memory_cell
X891 bl27 wl27 pl27 gnd memory_cell
X892 bl27 wl28 pl28 gnd memory_cell
X893 bl27 wl29 pl29 gnd memory_cell
X894 bl27 wl30 pl30 gnd memory_cell
X895 bl27 wl31 pl31 gnd memory_cell
X896 bl28 wl0 pl0 gnd memory_cell
X897 bl28 wl1 pl1 gnd memory_cell
X898 bl28 wl2 pl2 gnd memory_cell
X899 bl28 wl3 pl3 gnd memory_cell
X900 bl28 wl4 pl4 gnd memory_cell
X901 bl28 wl5 pl5 gnd memory_cell
X902 bl28 wl6 pl6 gnd memory_cell
X903 bl28 wl7 pl7 gnd memory_cell
X904 bl28 wl8 pl8 gnd memory_cell
X905 bl28 wl9 pl9 gnd memory_cell
X906 bl28 wl10 pl10 gnd memory_cell
X907 bl28 wl11 pl11 gnd memory_cell
X908 bl28 wl12 pl12 gnd memory_cell
X909 bl28 wl13 pl13 gnd memory_cell
X910 bl28 wl14 pl14 gnd memory_cell
X911 bl28 wl15 pl15 gnd memory_cell
X912 bl28 wl16 pl16 gnd memory_cell
X913 bl28 wl17 pl17 gnd memory_cell
X914 bl28 wl18 pl18 gnd memory_cell
X915 bl28 wl19 pl19 gnd memory_cell
X916 bl28 wl20 pl20 gnd memory_cell
X917 bl28 wl21 pl21 gnd memory_cell
X918 bl28 wl22 pl22 gnd memory_cell
X919 bl28 wl23 pl23 gnd memory_cell
X920 bl28 wl24 pl24 gnd memory_cell
X921 bl28 wl25 pl25 gnd memory_cell
X922 bl28 wl26 pl26 gnd memory_cell
X923 bl28 wl27 pl27 gnd memory_cell
X924 bl28 wl28 pl28 gnd memory_cell
X925 bl28 wl29 pl29 gnd memory_cell
X926 bl28 wl30 pl30 gnd memory_cell
X927 bl28 wl31 pl31 gnd memory_cell
X928 bl29 wl0 pl0 gnd memory_cell
X929 bl29 wl1 pl1 gnd memory_cell
X930 bl29 wl2 pl2 gnd memory_cell
X931 bl29 wl3 pl3 gnd memory_cell
X932 bl29 wl4 pl4 gnd memory_cell
X933 bl29 wl5 pl5 gnd memory_cell
X934 bl29 wl6 pl6 gnd memory_cell
X935 bl29 wl7 pl7 gnd memory_cell
X936 bl29 wl8 pl8 gnd memory_cell
X937 bl29 wl9 pl9 gnd memory_cell
X938 bl29 wl10 pl10 gnd memory_cell
X939 bl29 wl11 pl11 gnd memory_cell
X940 bl29 wl12 pl12 gnd memory_cell
X941 bl29 wl13 pl13 gnd memory_cell
X942 bl29 wl14 pl14 gnd memory_cell
X943 bl29 wl15 pl15 gnd memory_cell
X944 bl29 wl16 pl16 gnd memory_cell
X945 bl29 wl17 pl17 gnd memory_cell
X946 bl29 wl18 pl18 gnd memory_cell
X947 bl29 wl19 pl19 gnd memory_cell
X948 bl29 wl20 pl20 gnd memory_cell
X949 bl29 wl21 pl21 gnd memory_cell
X950 bl29 wl22 pl22 gnd memory_cell
X951 bl29 wl23 pl23 gnd memory_cell
X952 bl29 wl24 pl24 gnd memory_cell
X953 bl29 wl25 pl25 gnd memory_cell
X954 bl29 wl26 pl26 gnd memory_cell
X955 bl29 wl27 pl27 gnd memory_cell
X956 bl29 wl28 pl28 gnd memory_cell
X957 bl29 wl29 pl29 gnd memory_cell
X958 bl29 wl30 pl30 gnd memory_cell
X959 bl29 wl31 pl31 gnd memory_cell
X960 bl30 wl0 pl0 gnd memory_cell
X961 bl30 wl1 pl1 gnd memory_cell
X962 bl30 wl2 pl2 gnd memory_cell
X963 bl30 wl3 pl3 gnd memory_cell
X964 bl30 wl4 pl4 gnd memory_cell
X965 bl30 wl5 pl5 gnd memory_cell
X966 bl30 wl6 pl6 gnd memory_cell
X967 bl30 wl7 pl7 gnd memory_cell
X968 bl30 wl8 pl8 gnd memory_cell
X969 bl30 wl9 pl9 gnd memory_cell
X970 bl30 wl10 pl10 gnd memory_cell
X971 bl30 wl11 pl11 gnd memory_cell
X972 bl30 wl12 pl12 gnd memory_cell
X973 bl30 wl13 pl13 gnd memory_cell
X974 bl30 wl14 pl14 gnd memory_cell
X975 bl30 wl15 pl15 gnd memory_cell
X976 bl30 wl16 pl16 gnd memory_cell
X977 bl30 wl17 pl17 gnd memory_cell
X978 bl30 wl18 pl18 gnd memory_cell
X979 bl30 wl19 pl19 gnd memory_cell
X980 bl30 wl20 pl20 gnd memory_cell
X981 bl30 wl21 pl21 gnd memory_cell
X982 bl30 wl22 pl22 gnd memory_cell
X983 bl30 wl23 pl23 gnd memory_cell
X984 bl30 wl24 pl24 gnd memory_cell
X985 bl30 wl25 pl25 gnd memory_cell
X986 bl30 wl26 pl26 gnd memory_cell
X987 bl30 wl27 pl27 gnd memory_cell
X988 bl30 wl28 pl28 gnd memory_cell
X989 bl30 wl29 pl29 gnd memory_cell
X990 bl30 wl30 pl30 gnd memory_cell
X991 bl30 wl31 pl31 gnd memory_cell
X992 bl31 wl0 pl0 gnd memory_cell
X993 bl31 wl1 pl1 gnd memory_cell
X994 bl31 wl2 pl2 gnd memory_cell
X995 bl31 wl3 pl3 gnd memory_cell
X996 bl31 wl4 pl4 gnd memory_cell
X997 bl31 wl5 pl5 gnd memory_cell
X998 bl31 wl6 pl6 gnd memory_cell
X999 bl31 wl7 pl7 gnd memory_cell
X1000 bl31 wl8 pl8 gnd memory_cell
X1001 bl31 wl9 pl9 gnd memory_cell
X1002 bl31 wl10 pl10 gnd memory_cell
X1003 bl31 wl11 pl11 gnd memory_cell
X1004 bl31 wl12 pl12 gnd memory_cell
X1005 bl31 wl13 pl13 gnd memory_cell
X1006 bl31 wl14 pl14 gnd memory_cell
X1007 bl31 wl15 pl15 gnd memory_cell
X1008 bl31 wl16 pl16 gnd memory_cell
X1009 bl31 wl17 pl17 gnd memory_cell
X1010 bl31 wl18 pl18 gnd memory_cell
X1011 bl31 wl19 pl19 gnd memory_cell
X1012 bl31 wl20 pl20 gnd memory_cell
X1013 bl31 wl21 pl21 gnd memory_cell
X1014 bl31 wl22 pl22 gnd memory_cell
X1015 bl31 wl23 pl23 gnd memory_cell
X1016 bl31 wl24 pl24 gnd memory_cell
X1017 bl31 wl25 pl25 gnd memory_cell
X1018 bl31 wl26 pl26 gnd memory_cell
X1019 bl31 wl27 pl27 gnd memory_cell
X1020 bl31 wl28 pl28 gnd memory_cell
X1021 bl31 wl29 pl29 gnd memory_cell
X1022 bl31 wl30 pl30 gnd memory_cell
X1023 bl31 wl31 pl31 gnd memory_cell
X1024 bl0 ref seb nb nt vdd gnd sense_amp
X1025 bl1 ref seb nb nt vdd gnd sense_amp
X1026 bl2 ref seb nb nt vdd gnd sense_amp
X1027 bl3 ref seb nb nt vdd gnd sense_amp
X1028 bl4 ref seb nb nt vdd gnd sense_amp
X1029 bl5 ref seb nb nt vdd gnd sense_amp
X1030 bl6 ref seb nb nt vdd gnd sense_amp
X1031 bl7 ref seb nb nt vdd gnd sense_amp
X1032 bl8 ref seb nb nt vdd gnd sense_amp
X1033 bl9 ref seb nb nt vdd gnd sense_amp
X1034 bl10 ref seb nb nt vdd gnd sense_amp
X1035 bl11 ref seb nb nt vdd gnd sense_amp
X1036 bl12 ref seb nb nt vdd gnd sense_amp
X1037 bl13 ref seb nb nt vdd gnd sense_amp
X1038 bl14 ref seb nb nt vdd gnd sense_amp
X1039 bl15 ref seb nb nt vdd gnd sense_amp
X1040 bl16 ref seb nb nt vdd gnd sense_amp
X1041 bl17 ref seb nb nt vdd gnd sense_amp
X1042 bl18 ref seb nb nt vdd gnd sense_amp
X1043 bl19 ref seb nb nt vdd gnd sense_amp
X1044 bl20 ref seb nb nt vdd gnd sense_amp
X1045 bl21 ref seb nb nt vdd gnd sense_amp
X1046 bl22 ref seb nb nt vdd gnd sense_amp
X1047 bl23 ref seb nb nt vdd gnd sense_amp
X1048 bl24 ref seb nb nt vdd gnd sense_amp
X1049 bl25 ref seb nb nt vdd gnd sense_amp
X1050 bl26 ref seb nb nt vdd gnd sense_amp
X1051 bl27 ref seb nb nt vdd gnd sense_amp
X1052 bl28 ref seb nb nt vdd gnd sense_amp
X1053 bl29 ref seb nb nt vdd gnd sense_amp
X1054 bl30 ref seb nb nt vdd gnd sense_amp
X1055 bl31 ref seb nb nt vdd gnd sense_amp
X1056 bl0 in bl_gnd vdd gnd top_driver
X1057 bl1 in bl_gnd vdd gnd top_driver
X1058 bl2 in bl_gnd vdd gnd top_driver
X1059 bl3 in bl_gnd vdd gnd top_driver
X1060 bl4 in bl_gnd vdd gnd top_driver
X1061 bl5 in bl_gnd vdd gnd top_driver
X1062 bl6 in bl_gnd vdd gnd top_driver
X1063 bl7 in bl_gnd vdd gnd top_driver
X1064 bl8 in bl_gnd vdd gnd top_driver
X1065 bl9 in bl_gnd vdd gnd top_driver
X1066 bl10 in bl_gnd vdd gnd top_driver
X1067 bl11 in bl_gnd vdd gnd top_driver
X1068 bl12 in bl_gnd vdd gnd top_driver
X1069 bl13 in bl_gnd vdd gnd top_driver
X1070 bl14 in bl_gnd vdd gnd top_driver
X1071 bl15 in bl_gnd vdd gnd top_driver
X1072 bl16 in bl_gnd vdd gnd top_driver
X1073 bl17 in bl_gnd vdd gnd top_driver
X1074 bl18 in bl_gnd vdd gnd top_driver
X1075 bl19 in bl_gnd vdd gnd top_driver
X1076 bl20 in bl_gnd vdd gnd top_driver
X1077 bl21 in bl_gnd vdd gnd top_driver
X1078 bl22 in bl_gnd vdd gnd top_driver
X1079 bl23 in bl_gnd vdd gnd top_driver
X1080 bl24 in bl_gnd vdd gnd top_driver
X1081 bl25 in bl_gnd vdd gnd top_driver
X1082 bl26 in bl_gnd vdd gnd top_driver
X1083 bl27 in bl_gnd vdd gnd top_driver
X1084 bl28 in bl_gnd vdd gnd top_driver
X1085 bl29 in bl_gnd vdd gnd top_driver
X1086 bl30 in bl_gnd vdd gnd top_driver
X1087 bl31 in bl_gnd vdd gnd top_driver
* End of netlist. Compiled by NCS Memory compiler.