
* cell 
.SUBCKT 
.ENDS 
