# SA
.SUBCKT sense_amp in ref nt nb vdd gnd
.ENDS